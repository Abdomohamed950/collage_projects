library verilog;
use verilog.vl_types.all;
entity up_down_counter_dut is
end up_down_counter_dut;
