library verilog;
use verilog.vl_types.all;
entity testtt is
end testtt;
