library verilog;
use verilog.vl_types.all;
entity t_count_dut is
end t_count_dut;
