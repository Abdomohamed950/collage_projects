library verilog;
use verilog.vl_types.all;
entity test11 is
end test11;
